LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
LIBRARY WORK;

ENTITY MEMORYSTAGE_TEST IS   
	PORT( 
		-- INPUTS FROM MAIN MODULE
     	M_CLK : IN STD_LOGIC;
        M_RST : IN STD_LOGIC;
        M_INTERRUPT : IN STD_LOGIC;
        
        M_FETCHPC : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
        M_EXECUTEPC : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
        M_SIGNEXTENT : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
        M_ALURESULT : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
        
        M_MEMORYSIGNALS : IN STD_LOGIC_VECTOR (3 DOWNTO 0); -- 1 READ -- 1 WRITE -- 2 MUX SELECTOR
        M_PCORALU : IN STD_LOGIC; 
        M_GROUP1SELECTOR : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
        M_GROUP2SELECTOR : IN STD_LOGIC;  
        M_FLAGREGISTERIN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
        
        -- OUTPUTS TO MAIN MODULE
        M_FLAGREGISTEROUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        M_NEWFLAGDONE : OUT STD_LOGIC;
        M_NEWPC : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
        M_NEWPCDONE : OUT STD_LOGIC;
        M_MEMORYSTAGERESULT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
  
END ENTITY MEMORYSTAGE_TEST; 

ARCHITECTURE TESTARCH OF MEMORYSTAGE_TEST IS
  -- put declarations here.   
  -- INPUTS FROM DATAMEMORY MODULE
     SIGNAL S_DATAMEMORYDONEREAD : STD_LOGIC;
     SIGNAL S_DATAMEMORYDONEWRITE : STD_LOGIC;
     SIGNAL S_DATAMEMORYDATAOUT : STD_LOGIC_VECTOR (31 DOWNTO 0);  
     
     
        -- OUTPUTS TO DATAMEMORY MODULE
     SIGNAL S_DATAMEMORYREAD : STD_LOGIC;
     SIGNAL S_DATAMEMORYWRITE : STD_LOGIC;
     SIGNAL S_DATAMEMORYADDRESS : STD_LOGIC_VECTOR (10 DOWNTO 0); -- 
     SIGNAL S_DATAMEMORYDATAIN : STD_LOGIC_VECTOR (31 DOWNTO 0);
  
  
BEGIN
  -- put concurrent statements here.       
  MEMORY : ENTITY WORK.MEMORYMODULE generic map(32) port map (M_CLK,S_DATAMEMORYREAD, S_DATAMEMORYWRITE, S_DATAMEMORYDATAIN
                                    , S_DATAMEMORYADDRESS, S_DATAMEMORYDONEREAD, S_DATAMEMORYDONEWRITE, S_DATAMEMORYDATAOUT );
  
  MEMORYSTAGE : ENTITY WORK.MEMORY_STAGE  port map (M_CLK, M_RST, M_INTERRUPT, M_FETCHPC, M_EXECUTEPC, M_SIGNEXTENT, M_ALURESULT,
        							M_MEMORYSIGNALS, M_PCORALU, M_GROUP1SELECTOR, M_GROUP2SELECTOR,M_FLAGREGISTERIN,  S_DATAMEMORYDONEREAD,
        							S_DATAMEMORYDONEWRITE, S_DATAMEMORYDATAOUT, S_DATAMEMORYREAD, S_DATAMEMORYWRITE,
        							S_DATAMEMORYADDRESS,S_DATAMEMORYDATAIN,
        							M_FLAGREGISTEROUT, M_NEWFLAGDONE, M_NEWPC , M_NEWPCDONE, M_MEMORYSTAGERESULT );
        
  
END ARCHITECTURE TESTARCH; -- Of entity MEMORYSTAGE_TEST


