LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
LIBRARY WORK;

ENTITY MEMORYMODULE IS 
	GENERIC (DATASIZE : INTEGER := 16);
    PORT (
    	-- INPUTS
    	M_CLK : IN STD_LOGIC;
        M_READ : IN STD_LOGIC;
        M_WRITE : IN STD_LOGIC;
    	M_DATAIN : IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
        M_ADDRESS : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
        -- OUTPUTS
	    M_DONEREAD : OUT STD_LOGIC;
	    M_DONEWRITE : OUT STD_LOGIC;
        M_DATAOUT : OUT STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0)
        
    );
END ENTITY;

ARCHITECTURE MEMORYMODULEARCH OF MEMORYMODULE IS 

	 -- INPUT SIGNALS TO RAM  
      SIGNAL RAM_CLK : STD_LOGIC;
      SIGNAL RAM_MEMREAD : STD_LOGIC;
      SIGNAL RAM_MEMWRITE :  STD_LOGIC;
      SIGNAL RAM_ADDRESS : STD_LOGIC_VECTOR(11-1 DOWNTO 0);
      SIGNAL RAM_DATAIN :  STD_LOGIC_VECTOR(127 DOWNTO 0);
      
      -- OUTPUT SIGNALS FROM RAM 
      SIGNAL RAM_DATAOUT : STD_LOGIC_VECTOR(127 DOWNTO 0);
      SIGNAL RAM_READYSIGNAL :  STD_LOGIC;
      SIGNAL RAM_DONEWRITING :  STD_LOGIC;
      
      -- INPUT SIGNALS TO CACHE
  	  SIGNAL CACHE_CLK : STD_LOGIC;
      SIGNAL CACHE_INDEX :  STD_LOGIC_VECTOR (4 DOWNTO 0);
      SIGNAL CACHE_DISPLACEMENT : STD_LOGIC_VECTOR (2 DOWNTO 0);
      SIGNAL CACHE_CONTROLLERDATAIN :  STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
      SIGNAL CACHE_RAMDATAIN :  STD_LOGIC_VECTOR (127 DOWNTO 0);
      SIGNAL CACHE_CACHEREAD : STD_LOGIC;
      SIGNAL CACHE_CACHEWRITE : STD_LOGIC;
      SIGNAL CACHE_MEMORYREAD : STD_LOGIC;
      SIGNAL CACHE_MEMORYWRITE : STD_LOGIC;
      
      -- OUTPUT SIGNALS FROM CACHE
      SIGNAL CACHE_DATAOUT : STD_LOGIC_VECTOR(DATASIZE-1 DOWNTO 0);
      SIGNAL CACHE_MEMORYOUT : STD_LOGIC_VECTOR (127 DOWNTO 0);
      SIGNAL CACHE_DONEMEMORYREAD : STD_LOGIC;
      SIGNAL CACHE_DONEMEMORYWRITE : STD_LOGIC;
      SIGNAL CACHE_DONEREADSIGNAL : STD_LOGIC;
      SIGNAL CACHE_DONEWRITESIGNAL : STD_LOGIC;
      
       -- INPUT SIGNALS TO CONTROLLER 
  	SIGNAL CONTROLLER_CLK : STD_LOGIC;
    SIGNAL CONTROLLER_ADDRESSIN :  STD_LOGIC_VECTOR (10 DOWNTO 0);
    SIGNAL CONTROLLER_DATAIN :   STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
    SIGNAL CONTROLLER_READSIGNAL :  STD_LOGIC;
    SIGNAL CONTROLLER_WRITESIGNAL :  STD_LOGIC;
    SIGNAL CONTROLLER_MEMORYREADY :  STD_LOGIC;
    SIGNAL CONTROLLER_MEMORYDONEWRITING :  STD_LOGIC;
    SIGNAL CONTROLLER_CACHEDONEMEMORYREAD : STD_LOGIC;
    SIGNAL CONTROLLER_CACHEDONEMEMORYWRITE : STD_LOGIC;
    -- OUTPUT SIGNALS FROM CONTROLLER
    SIGNAL CONTROLLER_MEMREAD :  STD_LOGIC;
    SIGNAL CONTROLLER_MEMWRITE :  STD_LOGIC;
    SIGNAL CONTROLLER_ADDRESSOUT :  STD_LOGIC_VECTOR (10 DOWNTO 0);
    SIGNAL CONTROLLER_CACHEREAD :  STD_LOGIC;
    SIGNAL CONTROLLER_CACHEWRITE :  STD_LOGIC;
    SIGNAL CONTROLLER_CACHETOMEMWRITE :  STD_LOGIC;
    SIGNAL CONTROLLER_CACHEFROMMEMREAD :  STD_LOGIC;
    SIGNAL CONTROLLER_INDEX :  STD_LOGIC_VECTOR (4 DOWNTO 0);
    SIGNAL CONTROLLER_DISPLACEMENT :  STD_LOGIC_VECTOR (2 DOWNTO 0 );
    SIGNAL CONTROLLER_CONTROLLERDATAOUT :  STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);   

	BEGIN
    CONTROLLER_U : ENTITY WORK.CACHECONTROLLER GENERIC MAP (DATASIZE) PORT MAP (CONTROLLER_CLK, CONTROLLER_ADDRESSIN, CONTROLLER_DATAIN, CONTROLLER_READSIGNAL, CONTROLLER_WRITESIGNAL, CONTROLLER_MEMORYREADY,CONTROLLER_MEMORYDONEWRITING, CONTROLLER_CACHEDONEMEMORYREAD, CONTROLLER_CACHEDONEMEMORYWRITE, CONTROLLER_MEMREAD, CONTROLLER_MEMWRITE,CONTROLLER_ADDRESSOUT, CONTROLLER_CACHEREAD, CONTROLLER_CACHEWRITE, CONTROLLER_CACHETOMEMWRITE, CONTROLLER_CACHEFROMMEMREAD, CONTROLLER_INDEX, CONTROLLER_DISPLACEMENT, CONTROLLER_CONTROLLERDATAOUT );

    CACHE_U : ENTITY WORK.CACHE GENERIC MAP (DATASIZE) PORT MAP (CACHE_CLK, CACHE_INDEX, CACHE_DISPLACEMENT, CACHE_CONTROLLERDATAIN, CACHE_RAMDATAIN, CACHE_CACHEREAD, CACHE_CACHEWRITE,CACHE_MEMORYREAD, CACHE_MEMORYWRITE, CACHE_DATAOUT, CACHE_MEMORYOUT, CACHE_DONEMEMORYREAD, CACHE_DONEMEMORYWRITE, CACHE_DONEREADSIGNAL, CACHE_DONEWRITESIGNAL );
    
    RAM_U : ENTITY WORK.RAM PORT MAP (RAM_CLK, RAM_MEMREAD, RAM_MEMWRITE, RAM_ADDRESS, RAM_DATAIN,  RAM_DATAOUT, RAM_READYSIGNAL,RAM_DONEWRITING );
    
    PROCESS (M_CLK) IS
	BEGIN
    
    	  -- ASSIGNING CLOCKS TO EACH MODULE
          CONTROLLER_CLK <= M_CLK;
          CACHE_CLK <= M_CLK;
          RAM_CLK <= M_CLK;
          
          -- ASSIGNING CONTROLLER INPUT SIGNALS FROM MAIN MODULE
          CONTROLLER_ADDRESSIN <= M_ADDRESS;
          CONTROLLER_DATAIN <= M_DATAIN;
          CONTROLLER_READSIGNAL <= M_READ;
          CONTROLLER_WRITESIGNAL <= M_WRITE;
          
          -- ASSIGNING CACHE INPUT SIGNALS
          CACHE_INDEX <= CONTROLLER_INDEX ;
          CACHE_DISPLACEMENT <= CONTROLLER_DISPLACEMENT;
          CACHE_CONTROLLERDATAIN <= CONTROLLER_CONTROLLERDATAOUT;
          CACHE_CACHEREAD <= CONTROLLER_CACHEREAD;
          CACHE_CACHEWRITE <= CONTROLLER_CACHEWRITE;
          CACHE_MEMORYREAD <= CONTROLLER_CACHEFROMMEMREAD;
          CACHE_MEMORYWRITE <= CONTROLLER_CACHETOMEMWRITE;
          
          -- ASSIGNING RAM INPUT SIGNALS
          RAM_MEMREAD <= CONTROLLER_MEMREAD ;
          RAM_MEMWRITE <= CONTROLLER_MEMWRITE ;
          RAM_ADDRESS <= CONTROLLER_ADDRESSOUT;
          
          -- FOLLOW ASSIGNING CONTROLLER INPUT SIGNALS
          CONTROLLER_MEMORYREADY <= RAM_READYSIGNAL;
          CONTROLLER_MEMORYDONEWRITING <= RAM_DONEWRITING;
          CONTROLLER_CACHEDONEMEMORYREAD <= CACHE_DONEREADSIGNAL;
          CONTROLLER_CACHEDONEMEMORYWRITE <= CACHE_DONEWRITESIGNAL;
          
          -- FOLLOW ASSIGNING CACHE INPUT SIGNALS
          CACHE_RAMDATAIN <= RAM_DATAOUT;
          
          -- FOLLOW ASSIGNING RAM INPUT SIGNALS
          RAM_DATAIN <= CACHE_MEMORYOUT;
          
          -- ASSIGNING OUTPUTS OF MEMORYMODULE
          M_DONEREAD <= CACHE_DONEREADSIGNAL;
          M_DONEWRITE <= CACHE_DONEWRITESIGNAL;
          M_DATAOUT <= CACHE_DATAOUT;
    
    END PROCESS;



END MEMORYMODULEARCH;