LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY MEMORYMODULE IS 
	GENERIC (DATASIZE : INTEGER := 16);
    PORT (
    	M_CLK : IN STD_LOGIC;
        M_READ : IN STD_LOGIC;
        M_WRITE : IN STD_LOGIC;
    	M_DATAIN : IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
        M_ADDRESS : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
	M_DONEREAD : OUT STD_LOGIC;
        M_DATAOUT : OUT STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0)
        
    );
END ENTITY;

ARCHITECTURE MEMORYMODULEARCH OF MEMORYMODULE IS 
	
   

	COMPONENT CACHECONTROLLER IS 
      GENERIC (DATASIZE : INTEGER := 16);
      PORT (
        CLK : IN STD_LOGIC;
        ADDRESSIN : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
        DATAIN :  IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
        READSIGNAL : IN STD_LOGIC;
        WRITESIGNAL : IN STD_LOGIC;
        MEMREAD : OUT STD_LOGIC;
        MEMWRITE : OUT STD_LOGIC;
        CACHEREAD : OUT STD_LOGIC;
        CACHEWRITE : OUT STD_LOGIC;
        CACHETOMEMWRITE : OUT STD_LOGIC;
        ADDRESSOUT : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
        INDEX : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
        DISPLACEMENT : OUT STD_LOGIC_VECTOR (2 DOWNTO 0 );
        CONTROLLERDATAOUT : OUT STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0)

   	 );
    END COMPONENT CACHECONTROLLER;
    
    COMPONENT CACHE IS 
      GENERIC (DATASIZE : INTEGER := 16);
      PORT( 
          CLK : IN STD_LOGIC;
          INDEX : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
          DISPLACEMENT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
          CONTROLLERDATAIN : IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
          RAMDATAIN : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
          CACHEREAD : IN STD_LOGIC;
          CACHEWRITE : IN STD_LOGIC;
          MEMORYWRITE : IN STD_LOGIC;
          READYSIGNAL : IN STD_LOGIC;
	  DONESIGNAL : OUT STD_LOGIC;
          MEMORYOUT : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
          DATAOUT : OUT STD_LOGIC_VECTOR(DATASIZE-1 DOWNTO 0)
      );
    END COMPONENT CACHE;
    
    COMPONENT RAM IS
      GENERIC (ADDRESSWIDTH : INTEGER := 11; 
               RAMWIDTH : INTEGER := 16;
               RAMHEIGHT : INTEGER := 2048);
      PORT(
        CLK : IN STD_LOGIC;
        MEMREAD : IN STD_LOGIC;
        MEMWRITE : IN STD_LOGIC;
        ADDRESS : IN STD_LOGIC_VECTOR(ADDRESSWIDTH-1 DOWNTO 0);
        DATAIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
        DATAOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
        READYSIGNAL : OUT STD_LOGIC
      );
    END COMPONENT RAM;
    
    -- OUT SIGNALS FOR CONTROLLER
    SIGNAL MEMORY_READ_SIGNAL, MEMORY_WRITE_SIGNAL, CACHE_READ_SIGNAL, CACHE_WRITE_SIGNAL, CACHE_TOMEM_WRITE_SIGNAL : STD_LOGIC := '0';
    SIGNAL CONTROLLER_ADDRESSOUT : STD_LOGIC_VECTOR (10 DOWNTO 0);
    SIGNAL CONTROLLER_INDEX_OUT : STD_LOGIC_VECTOR (4 DOWNTO 0);
    SIGNAL CONTROLLER_DISPLACEMENT_OUT : STD_LOGIC_VECTOR (2 DOWNTO 0);
    SIGNAL CONTROLLER_DATAOUT : STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
    
    -- OUT SIGNALS FOR CACHE
    SIGNAL CACHE_DONESIGNAL : STD_LOGIC;
    SIGNAL CACHE_MEMORYOUT :  STD_LOGIC_VECTOR (127 DOWNTO 0);
    SIGNAL CACHE_DATAOUT : STD_LOGIC_VECTOR(DATASIZE-1 DOWNTO 0);
    
    -- OUT SIGNALS FOR RAM
    SIGNAL RAM_DATAOUT : STD_LOGIC_VECTOR (127 DOWNTO 0);
    SIGNAL RAM_READYSIGNAL : STD_LOGIC;
    
	
    
  BEGIN
  
    M_DATAOUT <= CACHE_DATAOUT;
    M_DONEREAD <= CACHE_DONESIGNAL;

    CONTROLLER_U : CACHECONTROLLER GENERIC MAP (DATASIZE) PORT MAP (M_CLK, M_ADDRESS, M_DATAIN, M_READ, M_WRITE, MEMORY_READ_SIGNAL, MEMORY_WRITE_SIGNAL, CACHE_READ_SIGNAL, CACHE_WRITE_SIGNAL, CACHE_TOMEM_WRITE_SIGNAL, CONTROLLER_ADDRESSOUT, CONTROLLER_INDEX_OUT, CONTROLLER_DISPLACEMENT_OUT, CONTROLLER_DATAOUT);

    CACHE_U : CACHE GENERIC MAP (DATASIZE) PORT MAP (M_CLK, CONTROLLER_INDEX_OUT, CONTROLLER_DISPLACEMENT_OUT, CONTROLLER_DATAOUT, RAM_DATAOUT, CACHE_READ_SIGNAL, CACHE_WRITE_SIGNAL, CACHE_TOMEM_WRITE_SIGNAL, RAM_READYSIGNAL, CACHE_DONESIGNAL, CACHE_MEMORYOUT, CACHE_DATAOUT );
    
    RAM_U : RAM GENERIC MAP (11, 16, 2048) PORT MAP (M_CLK, MEMORY_READ_SIGNAL, MEMORY_WRITE_SIGNAL, M_ADDRESS, CACHE_MEMORYOUT, RAM_DATAOUT );


END MEMORYMODULEARCH;