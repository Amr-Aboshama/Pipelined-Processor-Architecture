
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY CACHECONTROLLER IS 
  GENERIC (DATASIZE : INTEGER := 16);
  PORT (
    CLK : IN STD_LOGIC;
    ADDRESSIN : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
    DATAIN :  IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
    READSIGNAL : IN STD_LOGIC;
    WRITESIGNAL : IN STD_LOGIC;
    MEMREAD : OUT STD_LOGIC;
    MEMWRITE : OUT STD_LOGIC;
    CACHEREAD : OUT STD_LOGIC;
    CACHEWRITE : OUT STD_LOGIC;
    CACHETOMEMWRITE : OUT STD_LOGIC;
    ADDRESSOUT : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    INDEX : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    DISPLACEMENT : OUT STD_LOGIC_VECTOR (2 DOWNTO 0 );
    CONTROLLERDATAOUT : OUT STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0)

);
END ENTITY CACHECONTROLLER;

ARCHITECTURE CONTROLLERARCH OF CACHECONTROLLER IS 

  TYPE TAGSTYPE IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR (2 DOWNTO 0);
  TYPE DISPLACEMENTTYPE IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL TAGS : TAGSTYPE;
  SIGNAL DISP : DISPLACEMENTTYPE;
  SIGNAL VALID : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL DIRTY: STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL WRITESELFLATCH : STD_LOGIC := '0';
  SIGNAL READSELFLATCH : STD_LOGIC := '0';
  SIGNAL COUNTERWRITE0 : INTEGER RANGE 0 TO 5 := 0;
  SIGNAL COUNTERWRITE1 : INTEGER RANGE 0 TO 9 := 0;
  SIGNAL COUNTERREAD0 : INTEGER RANGE 0 TO 5 :=0;
  SIGNAL COUNTERREAD1 : INTEGER RANGE 0 TO 5 :=0;
  SIGNAL ADDRESSBUFFER : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL DATAINBUFFER : STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
  SIGNAL DIRTYTRIGGER1 : STD_LOGIC := '0';
  SIGNAL DIRTYTRIGGER2 : STD_LOGIC := '0';

  BEGIN

  PROCESS (CLK) IS
  
    BEGIN
    IF ( FALLING_EDGE(CLK)) THEN
      CACHEREAD <= '0';
      CACHEWRITE <= '0';
      MEMREAD <= '0';
      MEMWRITE <= '0';
      CACHETOMEMWRITE <= '0';
      IF (READSIGNAL = '1' OR WRITESIGNAL = '1') THEN
        ADDRESSBUFFER <= ADDRESSIN;
        DATAINBUFFER <= DATAIN;
      END IF;



      -- WRITE AND HIT
      IF (WRITESIGNAL = '1' AND VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) = '1' AND TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) = ADDRESSBUFFER(10 DOWNTO 8) ) THEN
        INDEX <= ADDRESSBUFFER(7 DOWNTO 3);
        DISPLACEMENT <= ADDRESSBUFFER(2 DOWNTO 0);
        CONTROLLERDATAOUT <= DATAINBUFFER;
        CACHEWRITE <= '1';
        DISP(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= ADDRESSBUFFER(2 DOWNTO 0);
      	DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= '1';
        VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= '1';

      -- WRITE AND MISS 
      ELSIF ((WRITESIGNAL = '1' OR WRITESELFLATCH = '1') AND (VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) /= '1' OR TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) /= ADDRESSBUFFER(10 DOWNTO 8))) THEN
     
        IF (DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) = '1' AND DIRTYTRIGGER2 = '0') THEN
            IF(COUNTERWRITE0 = 0) THEN -- FIRST MEMORY CYCLE (CACHE TO MEMORY)
                MEMWRITE <= '1';
                ADDRESSOUT <= TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) & ADDRESSBUFFER(7 DOWNTO 3) & "000";
                CACHETOMEMWRITE <= '1';
                INDEX <= ADDRESSBUFFER(7 DOWNTO 3);
		WRITESELFLATCH <= '1';
                COUNTERWRITE0 <= COUNTERWRITE0 +1;
            ELSIF (COUNTERWRITE0 = 1) THEN -- SECOND MEMORY CYCLE (CACHE TO MEMORY)
                COUNTERWRITE0 <= COUNTERWRITE0 +1;
            ELSIF (COUNTERWRITE0 = 2) THEN -- THIRD MEMORY CYCLE (CACHE TO MEMORY)
                COUNTERWRITE0 <= COUNTERWRITE0 +1;
            ELSIF (COUNTERWRITE0 = 3) THEN -- FOURTH MEMORY CYCLE (CACHE TO MEMORY)
            	DIRTYTRIGGER2 <= '1';
                COUNTERWRITE0 <= COUNTERWRITE0 +1;
            END IF; -- IF FOR COUNTERWRITE0
            
        ELSIF (DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) /= '1' OR DIRTYTRIGGER2 = '1') THEN
            IF (COUNTERWRITE1 = 0) THEN  --FIRST MEM CYCLE (MEMORY TO CACHE)
              MEMREAD <= '1';
              ADDRESSOUT <= ADDRESSIN(10 DOWNTO 3) & "000";
              WRITESELFLATCH <= '1';
              COUNTERWRITE1 <= COUNTERWRITE1 +1;
            ELSIF ( COUNTERWRITE1 = 1) THEN --SECOND MEMORY CYCLE (MEMORY TO CACHE)
              COUNTERWRITE1 <= COUNTERWRITE1 +1;
            ELSIF ( COUNTERWRITE1 = 2) THEN -- THIRD MEMORY CYCLE (MEMORY TO CACHE)
              COUNTERWRITE1 <= COUNTERWRITE1 +1;
            ELSIF ( COUNTERWRITE1 = 3) THEN -- FOURTH MEMORY CYCLE (MEMORY TO CACHE)
              COUNTERWRITE1 <= COUNTERWRITE1 +1;
            ELSIF ( COUNTERWRITE1 = 4) THEN -- CACHE READS FROM MEMORY 128 BITS (1 BLOCK)
              COUNTERWRITE1 <= COUNTERWRITE1 +1;
            ELSIF ( COUNTERWRITE1 = 5) THEN -- WRITE INTO CACHE THE NEW DATAIN
              CACHEWRITE <= '1';
              CONTROLLERDATAOUT <= DATAINBUFFER;
              INDEX <= ADDRESSBUFFER(7 DOWNTO 3);
              DISPLACEMENT <= ADDRESSBUFFER(2 DOWNTO 0);
              TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= ADDRESSBUFFER(10 DOWNTO 8);
              DISP(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= ADDRESSBUFFER(2 DOWNTO 0);
              VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= '1';
              DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= '1';
              WRITESELFLATCH <= '0';
	      DIRTYTRIGGER2 <= '0';
              COUNTERWRITE1 <= 0;
            END IF; -- IF FOR COUNTERWRITE1
          
        END IF; -- CHECK ON DIRTY BIT 
      
      -- READ AND HIT
      ELSIF (READSIGNAL = '1' AND VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) = '1' AND TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) = ADDRESSBUFFER(10 DOWNTO 8) ) THEN 
        INDEX <= ADDRESSBUFFER(7 DOWNTO 3);
        DISPLACEMENT <= ADDRESSBUFFER(2 DOWNTO 0);
      	CACHEREAD <= '1';

      -- READ AND MISS
      ELSIF ((READSIGNAL = '1' OR READSELFLATCH = '1') AND (VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) /= '1' OR TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) /= ADDRESSBUFFER(10 DOWNTO 8) )) THEN 
        IF (DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) = '1' AND DIRTYTRIGGER1 = '0') THEN 
        	IF (COUNTERREAD0 = 0) THEN -- FIRST MEMORY CYCLE (CACHE TO MEMORY)
            	MEMWRITE <= '1';
                ADDRESSOUT <= TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) & ADDRESSBUFFER(7 DOWNTO 3) & "000";
                CACHETOMEMWRITE <= '1';
                INDEX <= ADDRESSBUFFER(7 DOWNTO 3);
		READSELFLATCH <= '1';
                COUNTERREAD0 <= COUNTERREAD0 +1;
           	ELSIF (COUNTERREAD0 = 1) THEN -- SECOND MEMORY CYCLE (CACHE TO MEMORY)
            	COUNTERREAD0 <= COUNTERREAD0 +1;
           	ELSIF (COUNTERREAD0 = 2) THEN -- SECOND MEMORY CYCLE (CACHE TO MEMORY)
            	COUNTERREAD0 <= COUNTERREAD0 +1;
          	ELSIF (COUNTERREAD0 = 3) THEN -- SECOND MEMORY CYCLE (CACHE TO MEMORY)
            	DIRTYTRIGGER1 <= '1';
            	COUNTERREAD0 <= 0;
		END IF; -- END IF COUNTERREAD0
        
        ELSIF (DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) /= '1' OR DIRTYTRIGGER1 = '1') THEN
          IF ( COUNTERREAD1 = 0) THEN -- FIRST MEMORY CYCLE (MEMORY TO CACHE)
              MEMREAD <= '1';
              ADDRESSOUT <= ADDRESSBUFFER(10 DOWNTO 3) & "000";
              COUNTERREAD1 <= COUNTERREAD1 +1;
              READSELFLATCH <= '1';
          ELSIF (COUNTERREAD1 = 1) THEN -- SECOND MEMORY CYCLE (MEMORY TO CACHE)
              COUNTERREAD1 <= COUNTERREAD1 +1;
          ELSIF (COUNTERREAD1 = 2) THEN -- THIRD MEMORY CYCLE (MEMORY TO CACHE)
              COUNTERREAD1 <= COUNTERREAD1 +1;
          ELSIF (COUNTERREAD1 = 3) THEN -- FOURTH MEMORY CYCLE (MEMORY TO CACHE)
              COUNTERREAD1 <= COUNTERREAD1 +1;
          ELSIF (COUNTERREAD1 = 4) THEN -- CACHE READS FROM MEMORY 128 BITS (A WHOLE BLOCK)
              COUNTERREAD1 <= COUNTERREAD1 +1;
          ELSIF (COUNTERREAD1 = 5) THEN -- LET THE CACHE OUTPUT THE REQUIRED DATA
          	  CACHEREAD <= '1';
              INDEX <= ADDRESSBUFFER(7 DOWNTO 3);
              DISPLACEMENT <= ADDRESSBUFFER(2 DOWNTO 0);
              TAGS(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= ADDRESSBUFFER(10 DOWNTO 8);
              DISP(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= ADDRESSBUFFER(2 DOWNTO 0);
              DIRTY(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= '0';
              VALID(TO_INTEGER(UNSIGNED(ADDRESSBUFFER(7 DOWNTO 3)))) <= '1';
              READSELFLATCH <= '0';
              DIRTYTRIGGER1 <= '0';
              COUNTERREAD1 <= 0;
          END IF; -- COUNTERREAD1 IF     
        END IF; -- IF INSIDE READ AND MISS  
         	
     END IF; -- END OF 4 CASES

    END IF; -- FALLING EDGE
  END PROCESS;

END CONTROLLERARCH;









