LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
use std.textio.all;

ENTITY RAM IS
    GENERIC(
        DATA_WIDTH: INTEGER := 16;
        ADDRESS_WIDTH:  INTEGER := 11
    );
    
	PORT (
      -- INPUTS 
      CLK : IN STD_LOGIC;
      MEMREAD : IN STD_LOGIC;
      MEMWRITE : IN STD_LOGIC;
      ADDRESS : IN STD_LOGIC_VECTOR(11-1 DOWNTO 0);
      DATAIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
      
      -- OUTPUTS 
      DATAOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
      READYSIGNAL : OUT STD_LOGIC;
      DONEWRITING : OUT STD_LOGIC
      
    );

END ENTITY;

ARCHITECTURE RAMARCH OF RAM IS 

	-- RAM ITSELF 
    TYPE MEMORYTYPE IS ARRAY ((2**ADDRESS_WIDTH)-1 DOWNTO 0) OF STD_LOGIC_VECTOR (DATA_WIDTH-1 DOWNTO 0);

    IMPURE FUNCTION INIT_RAM_BIN RETURN MEMORYTYPE IS
        FILE TEXT_FILE : TEXT OPEN READ_MODE IS "FILE.bin";    --FILE NAME HERE
        VARIABLE TEXT_LINE : LINE;
        VARIABLE RAM_CONTENT : MEMORYTYPE;
        VARIABLE BV : BIT_VECTOR(RAM_CONTENT(0)'RANGE);
      BEGIN
        FOR I IN 0 TO (2**ADDRESS_WIDTH) - 1 LOOP
            IF(NOT ENDFILE(TEXT_FILE)) THEN
                READLINE(TEXT_FILE, TEXT_LINE);
                READ(TEXT_LINE, BV);
                RAM_CONTENT(I) := TO_STDLOGICVECTOR(BV);
            ELSE
                RAM_CONTENT(I) := (OTHERS=>'0') ;
            END IF;
        END LOOP;
        RETURN RAM_CONTENT;
      END FUNCTION;



    SIGNAL MEMORY : MEMORYTYPE := INIT_RAM_BIN;
    SIGNAL COUNTERWRITE : INTEGER RANGE 0 TO 3 := 0;
  	SIGNAL COUNTERREAD : INTEGER RANGE 0 TO 3 := 0;
    SIGNAL R_LATCH,W_LATCH : STD_LOGIC := '0';
    SIGNAL INBUFFER : STD_LOGIC_VECTOR(127 DOWNTO 0);
    SIGNAL OUTBUFFER : STD_LOGIC_VECTOR(127 DOWNTO 0);
    

    BEGIN 
    PROCESS (CLK) IS
    
    	BEGIN        
    	IF (RISING_EDGE(CLK)) THEN
        
        	READYSIGNAL <= '0';
       		DONEWRITING <= '0';
        	
        	-- WRITE TO MEMORY
        	IF (MEMWRITE = '1' OR W_LATCH = '1') THEN
                  IF (COUNTERWRITE = 0)THEN
                      INBUFFER <= DATAIN;
                      COUNTERWRITE <= COUNTERWRITE +1;
                      W_LATCH <= '1';
                  ELSIF (COUNTERWRITE = 1) THEN
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))) <= INBUFFER(15 DOWNTO 0);
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+1) <= INBUFFER(31 DOWNTO 16);
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+2) <= INBUFFER(47 DOWNTO 32);
                      COUNTERWRITE <= COUNTERWRITE +1;
                  ELSIF (COUNTERWRITE = 2) THEN
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+3) <= INBUFFER(63 DOWNTO 48);
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+4) <= INBUFFER(79 DOWNTO 64);
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+5) <= INBUFFER(95 DOWNTO 80);
                      COUNTERWRITE <= COUNTERWRITE +1;
                  ELSE 
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+6) <= INBUFFER(111 DOWNTO 96);
                      MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+7) <= INBUFFER(127 DOWNTO 112);
                      DONEWRITING <= '1';
                      COUNTERWRITE <= 0;
                      W_LATCH <= '0';
                  END IF; -- COUNTERWRITE


            -- READ FROM MEMORY
            ELSIF (MEMREAD = '1' OR R_LATCH = '1') THEN
              IF (COUNTERREAD = 0) THEN
                  OUTBUFFER(15 DOWNTO 0) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)));
                  OUTBUFFER(31 DOWNTO 16) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+1);
                  OUTBUFFER(47 DOWNTO 32) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+2);
                  COUNTERREAD <= COUNTERREAD +1;
                  R_LATCH <= '1';
              ELSIF (COUNTERREAD = 1) THEN
                  OUTBUFFER(63 DOWNTO 48) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+3);
                  OUTBUFFER(79 DOWNTO 64) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+4);
                  OUTBUFFER(95 DOWNTO 80) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+5);
                  COUNTERREAD <= COUNTERREAD +1;
              ELSIF (COUNTERREAD = 2) THEN
                  OUTBUFFER(111 DOWNTO 96) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+6);
                  OUTBUFFER(127 DOWNTO 112) <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))+7);
                  COUNTERREAD <= COUNTERREAD +1;
              ELSE
                  DATAOUT <= OUTBUFFER;
                  READYSIGNAL <= '1';
                  COUNTERREAD <= 0;
                  R_LATCH <= '0';
              END IF; -- COUNTER READ 
              
            END IF; -- READ OR WRITE
        
        END IF; -- FALLING EDGE
    
    END PROCESS;

END RAMARCH;