LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

entity BRANCH_PREDECTION_UNIT is
    port (
        
    ) ;
end BRANCH_PREDECTION_UNIT;