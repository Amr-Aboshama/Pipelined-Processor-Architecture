LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY CACHE IS 
  GENERIC (DATASIZE : INTEGER := 16);
  PORT( 
      CLK : IN STD_LOGIC;
      INDEX : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      DISPLACEMENT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      CONTROLLERDATAIN : IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
      RAMDATAIN : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
      CACHEREAD : IN STD_LOGIC;
      CACHEWRITE : IN STD_LOGIC;
      MEMORYWRITE : IN STD_LOGIC;
      READYSIGNAL : IN STD_LOGIC;
      DONEREADSIGNAL : OUT STD_LOGIC;
      DONEWRITESIGNAL : OUT STD_LOGIC;
      MEMORYOUT : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
      DATAOUT : OUT STD_LOGIC_VECTOR(DATASIZE-1 DOWNTO 0)
  );
END ENTITY CACHE;

ARCHITECTURE CACHEARCH OF CACHE IS 
  TYPE CACHETYPE IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR(127 DOWNTO 0);
  SIGNAL CACHE_S : CACHETYPE;
  SIGNAL SIG_RIGHT_INDEX : INTEGER RANGE 0 TO 255; -- FOR CHECKING
  SIGNAL SIG_LEFT_INDEX : INTEGER RANGE 0 TO 255; -- FOR CHECKING

  BEGIN
  PROCESS (CLK) IS
 
    VARIABLE RIGHT_INDEX : INTEGER RANGE 0 TO 255; 
    VARIABLE LEFT_INDEX : INTEGER RANGE 0 TO 255;
    
    BEGIN
    IF (FALLING_EDGE(CLK)) THEN 
      DONEREADSIGNAL <= '0';
      DONEWRITESIGNAL <= '0';
      LEFT_INDEX := DATASIZE - 1 + (TO_INTEGER(UNSIGNED(DISPLACEMENT))*DATASIZE) ;
      IF (LEFT_INDEX-DATASIZE+1 = 0 ) THEN 
        RIGHT_INDEX := 0;
      ELSE 
        RIGHT_INDEX := LEFT_INDEX-DATASIZE+1;
      END IF;

    SIG_LEFT_INDEX <= LEFT_INDEX; -- FOR CHECKING
    SIG_RIGHT_INDEX <= RIGHT_INDEX; -- FOR CHECKING


    IF (CACHEREAD = '1') THEN 
   	  DATAOUT <= CACHE_S(TO_INTEGER(UNSIGNED(INDEX)))(LEFT_INDEX DOWNTO RIGHT_INDEX);
	  DONEREADSIGNAL <= '1';
    ELSIF (CACHEWRITE = '1') THEN 
  	  CACHE_S(TO_INTEGER(UNSIGNED(INDEX)))(LEFT_INDEX DOWNTO RIGHT_INDEX)<= CONTROLLERDATAIN;
	  DONEWRITESIGNAL <= '1';
    ELSIF (READYSIGNAL = '1') THEN 
  	  CACHE_S(TO_INTEGER(UNSIGNED(INDEX)))<= RAMDATAIN;
    ELSIF (MEMORYWRITE = '1') THEN 
	  MEMORYOUT <= CACHE_S(TO_INTEGER(UNSIGNED(INDEX)));
    ELSE 
  	  DATAOUT <= "ZZZZZZZZZZZZZZZZ";
    END IF;
  END IF;
  END PROCESS;
END CACHEARCH;

