LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY MEMORYMODULE IS 
	GENERIC (DATASIZE : INTEGER := 16);
    PORT (
    	M_CLK : IN STD_LOGIC;
        M_READ : IN STD_LOGIC;
        M_WRITE : IN STD_LOGIC;
    	M_DATAIN : IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
        M_ADDRESS : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
	    M_DONEREAD : OUT STD_LOGIC;
	    M_DONEWRITE : OUT STD_LOGIC;
        M_DATAOUT : OUT STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0)
        
    );
END ENTITY;

ARCHITECTURE MEMORYMODULEARCH OF MEMORYMODULE IS 
	
   

	COMPONENT CACHECONTROLLER IS 
      GENERIC (DATASIZE : INTEGER := 16);
      PORT (
        CLK : IN STD_LOGIC;
        ADDRESSIN : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
        DATAIN :  IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
        READSIGNAL : IN STD_LOGIC;
        WRITESIGNAL : IN STD_LOGIC;
        MEMREAD : OUT STD_LOGIC;
        MEMWRITE : OUT STD_LOGIC;
        CACHEREAD : OUT STD_LOGIC;
        CACHEWRITE : OUT STD_LOGIC;
        CACHETOMEMWRITE : OUT STD_LOGIC;
        ADDRESSOUT : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
        INDEX : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
        DISPLACEMENT : OUT STD_LOGIC_VECTOR (2 DOWNTO 0 );
        CONTROLLERDATAOUT : OUT STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0)

   	 );
    END COMPONENT CACHECONTROLLER;
    
    COMPONENT CACHE IS 
      GENERIC (DATASIZE : INTEGER := 16);
      PORT( 
          CLK : IN STD_LOGIC;
          INDEX : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
          DISPLACEMENT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
          CONTROLLERDATAIN : IN STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
          RAMDATAIN : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
          CACHEREAD : IN STD_LOGIC;
          CACHEWRITE : IN STD_LOGIC;
          MEMORYWRITE : IN STD_LOGIC;
          READYSIGNAL : IN STD_LOGIC;
	      DONEREADSIGNAL : OUT STD_LOGIC;
          DONEWRITESIGNAL : OUT STD_LOGIC;
          MEMORYOUT : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
          DATAOUT : OUT STD_LOGIC_VECTOR(DATASIZE-1 DOWNTO 0)
      );
    END COMPONENT CACHE;
    
    COMPONENT RAM IS
      GENERIC (ADDRESSWIDTH : INTEGER := 11; 
               RAMWIDTH : INTEGER := 16;
               RAMHEIGHT : INTEGER := 2048);
      PORT(
        CLK : IN STD_LOGIC;
        MEMREAD : IN STD_LOGIC;
        MEMWRITE : IN STD_LOGIC;
        ADDRESS : IN STD_LOGIC_VECTOR(ADDRESSWIDTH-1 DOWNTO 0);
        DATAIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
        DATAOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
        READYSIGNAL : OUT STD_LOGIC
      );
    END COMPONENT RAM;
    
    -- IN AND OUT SIGNALS FOR CONTROLLER
    SIGNAL CONTROLLER_CLK :  STD_LOGIC;
    SIGNAL CONTROLLER_ADDRESSIN : STD_LOGIC_VECTOR (10 DOWNTO 0);
    SIGNAL CONTROLLER_DATAIN :  STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
    SIGNAL CONTROLLER_READSIGNAL : STD_LOGIC;
    SIGNAL CONTROLLER_WRITESIGNAL : STD_LOGIC;
    
    SIGNAL MEMORY_READ_SIGNAL, MEMORY_WRITE_SIGNAL, CACHE_READ_SIGNAL, CACHE_WRITE_SIGNAL, CACHE_TOMEM_WRITE_SIGNAL : STD_LOGIC := '0';
    SIGNAL CONTROLLER_ADDRESSOUT : STD_LOGIC_VECTOR (10 DOWNTO 0);
    SIGNAL CONTROLLER_INDEX_OUT : STD_LOGIC_VECTOR (4 DOWNTO 0);
    SIGNAL CONTROLLER_DISPLACEMENT_OUT : STD_LOGIC_VECTOR (2 DOWNTO 0);
    SIGNAL CONTROLLER_DATAOUT : STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
    
    -- IN AND OUT SIGNALS FOR CACHE
     SIGNAL CACHE_CLK : STD_LOGIC;
     SIGNAL CACHE_INDEX :  STD_LOGIC_VECTOR (4 DOWNTO 0);
     SIGNAL CACHE_DISPLACEMENT :  STD_LOGIC_VECTOR (2 DOWNTO 0);
     SIGNAL CACHE_CONTROLLERDATAIN : STD_LOGIC_VECTOR (DATASIZE-1 DOWNTO 0);
     SIGNAL CACHE_RAMDATAIN :  STD_LOGIC_VECTOR (127 DOWNTO 0);
     SIGNAL CACHE_CACHEREAD :  STD_LOGIC;
     SIGNAL CACHE_CACHEWRITE : STD_LOGIC;
     SIGNAL CACHE_MEMORYWRITE : STD_LOGIC;
     SIGNAL CACHE_READYSIGNAL :  STD_LOGIC;
    
    SIGNAL CACHE_DONEREADSIGNAL : STD_LOGIC;
    SIGNAL CACHE_DONEWRITESIGNAL : STD_LOGIC;
    SIGNAL CACHE_MEMORYOUT :  STD_LOGIC_VECTOR (127 DOWNTO 0);
    SIGNAL CACHE_DATAOUT : STD_LOGIC_VECTOR(DATASIZE-1 DOWNTO 0);
    
    -- IN AND OUT SIGNALS FOR RAM
    SIGNAL RAM_CLK :  STD_LOGIC;
    SIGNAL RAM_MEMREAD :  STD_LOGIC;
    SIGNAL RAM_MEMWRITE :  STD_LOGIC;
    SIGNAL RAM_ADDRESS :  STD_LOGIC_VECTOR(10 DOWNTO 0);
    SIGNAL RAM_DATAIN : STD_LOGIC_VECTOR(127 DOWNTO 0);
    
    SIGNAL RAM_DATAOUT : STD_LOGIC_VECTOR (127 DOWNTO 0);
    SIGNAL RAM_READYSIGNAL : STD_LOGIC;
    
	
    
  BEGIN
  
    M_DATAOUT <= CACHE_DATAOUT;
    M_DONEREAD <= CACHE_DONEREADSIGNAL;
    M_DONEWRITE <= CACHE_DONEWRITESIGNAL;

    CONTROLLER_U : CACHECONTROLLER GENERIC MAP (DATASIZE) PORT MAP (CONTROLLER_CLK, CONTROLLER_ADDRESSIN, CONTROLLER_DATAIN, CONTROLLER_READSIGNAL, CONTROLLER_WRITESIGNAL, MEMORY_READ_SIGNAL, MEMORY_WRITE_SIGNAL, CACHE_READ_SIGNAL, CACHE_WRITE_SIGNAL, CACHE_TOMEM_WRITE_SIGNAL, CONTROLLER_ADDRESSOUT, CONTROLLER_INDEX_OUT, CONTROLLER_DISPLACEMENT_OUT, CONTROLLER_DATAOUT);

    CACHE_U : CACHE GENERIC MAP (DATASIZE) PORT MAP (CACHE_CLK, CACHE_INDEX, CACHE_DISPLACEMENT, CACHE_CONTROLLERDATAIN, CACHE_RAMDATAIN, CACHE_CACHEREAD, CACHE_CACHEWRITE, CACHE_MEMORYWRITE, CACHE_READYSIGNAL, CACHE_DONEREADSIGNAL, CACHE_DONEWRITESIGNAL, CACHE_MEMORYOUT, CACHE_DATAOUT  );
    
    RAM_U : RAM GENERIC MAP (11, 16, 2048) PORT MAP (RAM_CLK, RAM_MEMREAD, RAM_MEMWRITE, RAM_ADDRESS, RAM_DATAIN,  RAM_DATAOUT, RAM_READYSIGNAL );

    PROCESS (M_CLK) IS
	BEGIN
    	--IF (RISING_EDGE(M_CLK)) THEN
        
        
          -- ASSIGNING CLOCKS TO EACH MODULE
          CONTROLLER_CLK <= M_CLK;
          CACHE_CLK <= M_CLK;
          RAM_CLK <= M_CLK;
          
          -- ASSIGNING CONTROLLER INPUT SIGNALS
          CONTROLLER_ADDRESSIN <= M_ADDRESS;
          CONTROLLER_DATAIN <= M_DATAIN;
          CONTROLLER_READSIGNAL <= M_READ;
          CONTROLLER_WRITESIGNAL <= M_WRITE;
          
          -- ASSIGNING CACHE INPUT SIGNALS
          CACHE_INDEX <= CONTROLLER_INDEX_OUT;
          CACHE_DISPLACEMENT <= CONTROLLER_DISPLACEMENT_OUT;
          CACHE_CONTROLLERDATAIN <= CONTROLLER_DATAOUT;
          CACHE_CACHEREAD <= CACHE_READ_SIGNAL;
          CACHE_CACHEWRITE <= CACHE_WRITE_SIGNAL;
          CACHE_MEMORYWRITE <= CACHE_TOMEM_WRITE_SIGNAL;
          
          
          -- ASSIGNING RAM INPUT SIGNALS
          RAM_MEMREAD <= MEMORY_READ_SIGNAL;
          RAM_MEMWRITE <= MEMORY_READ_SIGNAL;
          RAM_ADDRESS <= CONTROLLER_ADDRESSOUT;
          RAM_DATAIN <= CACHE_MEMORYOUT;
          
          -- FOLLOW CACHE INPUT SIGNALS
          CACHE_RAMDATAIN <= RAM_DATAOUT;
          CACHE_READYSIGNAL <= RAM_READYSIGNAL;

          -- CHANGING THE OUTPUT

          M_DATAOUT <= CACHE_DATAOUT;
    	  M_DONEREAD <= CACHE_DONEREADSIGNAL;
    	  M_DONEWRITE <= CACHE_DONEWRITESIGNAL;
          
          
    	--END IF;
    END PROCESS;

END MEMORYMODULEARCH;